// File: src/processor.sv
// Module: processor
// Purpose: Top level module for the processor.

module processor (
    // TODO: Add ports here
);
    //TODO: Instantiate submodules here once done
endmodule